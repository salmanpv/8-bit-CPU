// Accumulator

module accumulator (
    input wire clk,
    input wire reset,
    input wire load,
    input wire [7:0] data_in,
    output reg [7:0] data_out
);

    always @(posedge clk or posedge reset) begin
        if (reset)
            data_out <= 8'b0;  // Reset accumulator to 0
        else if (load)
            data_out <= data_in;  // Load new data into accumulator
    end
endmodule
